/* 
INSTALL V:
cd ~/bin
git clone https://github.com/vlang/v
cd v
make
sudo ./v symlink

RUN FILE:
v run main.v
*/

module main

fn main() {
	// display hello world
	println('Hello World!')
}
