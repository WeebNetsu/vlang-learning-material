/* 
INIT PROJECT:
v init - if already inside a folder
v new project - to create a new folder
v new project web - for a website template

RUN PROJECT

v run
or
cd src
v run main.v (your file name)

v main.v will build an executable
*/

module main

fn main() {
	// display hello world
	println('Hello World!')
}
